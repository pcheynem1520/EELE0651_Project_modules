module reducer_unit (
    /* input signals */

    /* input buses */
    
    /* output signal */
    
    /* output buses */
    
);

    

endmodule
