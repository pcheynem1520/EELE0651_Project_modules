module lower_zero_extender (
    /* input signals */

    /* input buses */
    
    /* output signal */
    
    /* output buses */
    
);

    

endmodule
