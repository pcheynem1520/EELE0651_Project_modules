//=========================================================
// EELE 0651: Computer Organization
// Authors: PJ Cheyne-Miller, Brenden O'Donnell
// Date: 10 November 2021
// Description:
// 
// Based on the clock signals and intruction being executed,
// it controls the chip enable and write enable signals of
// the processor memory.
//=========================================================

//module memory_signal_generator (
    /* input signals */
    //input logic clk,    // clock signal

    /* input buses */

    /* output signal */

    /* output buses */
    
//);
    
//endmodule
